`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03.05.2023 18:22:00
// Design Name: 
// Module Name: ALU_8_bit_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ALU_8_bit_tb();
reg [7:0] A;
reg [7:0] B;
reg [1:0] S1;
reg [2:0] S2;
reg [3:0] S3;
wire [7:0] O;
ALU_8_bit alu1(.A(A),.B(B),.S1(S1),.S2(S2),.S3(S3),.O(O));
initial
begin
A=8'b00000111;
B=8'b00000100;
S1=1'b0;
S2=3'b000;
S3=4'b0000;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b0;
S2=3'b001;
S3=4'b0000;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b0;
S2=3'b010;
S3=4'b0000;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b0;
S2=3'b011;
S3=4'b0000;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b0000;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b0001;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b0010;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b0011;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b0100;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b0101;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b0110;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b0111;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b1000;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b1001;
#10
A=8'b00000111;
B=8'b00000100;
S1=1'b1;
S2=3'b001;
S3=4'b1100;
end
endmodule
